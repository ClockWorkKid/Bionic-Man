* D:\My Documents\Documents\Google Drive\Projects\3. Bionic man\pspice2\Instrumentation.sch

* Schematics Version 9.2
* Sun Dec 02 01:55:48 2018



** Analysis setup **
.tran 1ns .2s 0
.OP 


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "Instrumentation.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
